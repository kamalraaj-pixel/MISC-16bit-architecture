module ram_initial();
input [255:0] ram;
assign ram[0]<=0;
assign ram[1]<=0;
assign ram[2]<=0;
assign ram[3]<=0;
assign ram[4]<=0;
assign ram[5]<=0;
assign ram[6]<=0;
assign ram[7]<=0;
assign ram[8]<=0;
assign ram[9]<=0;
assign ram[10]<=0;
assign ram[11]<=0;
assign ram[12]<=0;
assign ram[13]<=0;
assign ram[14]<=0;
assign ram[15]<=0;
assign ram[16]<=0;
assign ram[17]<=0;
assign ram[18]<=0;
assign ram[19]<=0;
assign ram[20]<=0;
assign ram[21]<=0;
assign ram[22]<=0;
assign ram[23]<=0;
assign ram[24]<=0;
assign ram[25]<=0;
assign ram[26]<=0;
assign ram[27]<=0;
assign ram[28]<=0;
assign ram[29]<=0;
assign ram[30]<=0;
assign ram[31]<=0;
assign ram[32]<=0;
assign ram[33]<=0;
assign ram[34]<=0;
assign ram[35]<=0;
assign ram[36]<=0;
assign ram[37]<=0;
assign ram[38]<=0;
assign ram[39]<=0;
assign ram[40]<=0;
assign ram[41]<=0;
assign ram[42]<=0;
assign ram[43]<=0;
assign ram[44]<=0;
assign ram[45]<=0;
assign ram[46]<=0;
assign ram[47]<=0;

assign ram[48]<=0;
assign ram[49]<=0;
assign ram[50]<=0;
assign ram[51]<=0;
assign ram[52]<=0;
assign ram[53]<=0;
assign ram[54]<=0;
assign ram[55]<=0;
assign ram[56]<=0;
assign ram[57]<=0;
assign ram[58]<=0;
assign ram[59]<=0;
assign ram[60]<=0;
assign ram[61]<=0;
assign ram[62]<=0;
assign ram[63]<=0;

assign ram[64]<=0;
assign ram[65]<=0;
assign ram[66]<=0;
assign ram[67]<=0;
assign ram[68]<=0;
assign ram[69]<=0;
assign ram[70]<=0;
assign ram[71]<=0;
assign ram[72]<=0;
assign ram[73]<=0;
assign ram[74]<=0;
assign ram[75]<=0;
assign ram[76]<=0;
assign ram[77]<=0;
assign ram[78]<=0;
assign ram[79]<=0;

assign ram[80]<=0;
assign ram[81]<=0;
assign ram[82]<=0;
assign ram[83]<=0;
assign ram[84]<=0;
assign ram[85]<=0;
assign ram[86]<=0;
assign ram[87]<=0;
assign ram[88]<=0;
assign ram[89]<=0;
assign ram[90]<=0;
assign ram[91]<=0;
assign ram[92]<=0;
assign ram[93]<=0;
assign ram[94]<=0;
assign ram[95]<=0;
assign ram[96]<=0;
assign ram[97]<=0;
assign ram[98]<=0;
assign ram[99]<=0;
assign ram[100]<=0;
assign ram[101]<=0;
assign ram[102]<=0;
assign ram[103]<=0;
assign ram[104]<=0;
assign ram[105]<=0;
assign ram[106]<=0;
assign ram[107]<=0;
assign ram[108]<=0;
assign ram[109]<=0;
assign ram[110]<=0;
assign ram[111]<=0;

assign ram[112]<=0;
assign ram[113]<=0;
assign ram[114]<=0;
assign ram[115]<=0;
assign ram[116]<=0;
assign ram[117]<=0;
assign ram[118]<=0;
assign ram[119]<=0;
assign ram[120]<=0;
assign ram[121]<=0;
assign ram[122]<=0;
assign ram[123]<=0;
assign ram[124]<=0;
assign ram[125]<=0;
assign ram[126]<=0;
assign ram[127]<=0;

assign ram[128]<=0;
assign ram[129]<=0;
assign ram[130]<=0;
assign ram[131]<=0;
assign ram[132]<=0;
assign ram[133]<=0;
assign ram[134]<=0;
assign ram[135]<=0;
assign ram[136]<=0;
assign ram[137]<=0;
assign ram[138]<=0;
assign ram[139]<=0;
assign ram[140]<=0;
assign ram[141]<=0;
assign ram[142]<=0;
assign ram[143]<=0;

assign ram[144]<=0;
assign ram[145]<=0;
assign ram[146]<=0;
assign ram[147]<=0;
assign ram[148]<=0;
assign ram[149]<=0;
assign ram[150]<=0;
assign ram[151]<=0;
assign ram[152]<=0;
assign ram[153]<=0;
assign ram[154]<=0;
assign ram[155]<=0;
assign ram[156]<=0;
assign ram[157]<=0;
assign ram[158]<=0;
assign ram[159]<=0;

assign ram[160]<=0;
assign ram[161]<=0;
assign ram[162]<=0;
assign ram[163]<=0;
assign ram[164]<=0;
assign ram[165]<=0;
assign ram[166]<=0;
assign ram[167]<=0;
assign ram[168]<=0;
assign ram[169]<=0;
assign ram[170]<=0;
assign ram[171]<=0;
assign ram[172]<=0;
assign ram[173]<=0;
assign ram[174]<=0;
assign ram[175]<=0;

assign ram[176]<=0;
assign ram[177]<=0;
assign ram[178]<=0;
assign ram[179]<=0;
assign ram[180]<=0;
assign ram[181]<=0;
assign ram[182]<=0;
assign ram[183]<=0;
assign ram[184]<=0;
assign ram[185]<=0;
assign ram[186]<=0;
assign ram[187]<=0;
assign ram[188]<=0;
assign ram[189]<=0;
assign ram[190]<=0;
assign ram[191]<=0;

assign ram[192]<=0;
assign ram[193]<=0;
assign ram[194]<=0;
assign ram[195]<=0;
assign ram[196]<=0;
assign ram[197]<=0;
assign ram[198]<=0;
assign ram[199]<=0;
assign ram[200]<=0;
assign ram[201]<=0;
assign ram[202]<=0;
assign ram[203]<=0;
assign ram[204]<=0;
assign ram[205]<=0;
assign ram[206]<=0;
assign ram[207]<=0;

assign ram[208]<=0;
assign ram[209]<=0;
assign ram[210]<=0;
assign ram[211]<=0;
assign ram[212]<=0;
assign ram[213]<=0;
assign ram[214]<=0;
assign ram[215]<=0;
assign ram[216]<=0;
assign ram[217]<=0;
assign ram[218]<=0;
assign ram[219]<=0;
assign ram[220]<=0;
assign ram[221]<=0;
assign ram[222]<=0;
assign ram[223]<=0;

assign ram[224]<=0;
assign ram[225]<=0;
assign ram[226]<=0;
assign ram[227]<=0;
assign ram[228]<=0;
assign ram[229]<=0;
assign ram[230]<=0;
assign ram[231]<=0;
assign ram[232]<=0;
assign ram[233]<=0;
assign ram[234]<=0;
assign ram[235]<=0;
assign ram[236]<=0;
assign ram[237]<=0;
assign ram[238]<=0;
assign ram[239]<=0;

assign ram[240]<=0;
assign ram[241]<=0;
assign ram[242]<=0;
assign ram[243]<=0;
assign ram[244]<=0;
assign ram[245]<=0;
assign ram[246]<=0;
assign ram[247]<=0;
assign ram[248]<=0;
assign ram[249]<=0;
assign ram[250]<=0;
assign ram[251]<=0;
assign ram[252]<=0;
assign ram[253]<=0;
assign ram[254]<=0;
assign ram[255]<=0;
end module




